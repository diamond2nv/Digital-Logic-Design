`timescale 1ns / 1ps


module myAND(
    input a,
    input b,
    output out
    );
    
    and g1(out,a,b);
endmodule
